`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Design Name: RISCV CPU
// Module Name: InstructionRamWrapper
// Target Devices: Nexys4
// Tool Versions: Vivado 2017.4.1
// Description: a Verilog-based ram which can be systhesis as BRAM
//////////////////////////////////////////////////////////////////////////////////
module InstructionRam(
    input  clk,
    input  web,
    input  [31:2] addra, addrb,
    input  [31:0] dinb,
    output reg [31:0] douta, doutb
);
initial begin douta=0; doutb=0; end

wire addra_valid = ( addra[31:14]==18'h0 );
wire addrb_valid = ( addrb[31:14]==18'h0 );
wire [11:0] addral = addra[13:2];
wire [11:0] addrbl = addrb[13:2];

reg [31:0] ram_cell [0:4095];

initial begin    // you can add simulation instructions here
    ram_cell[0] = 32'h00000000;
        // ......
end

always @ (posedge clk)
    douta <= addra_valid ? ram_cell[addral] : 0;
    
always @ (posedge clk)
    doutb <= addrb_valid ? ram_cell[addrbl] : 0;

always @ (posedge clk)
    if(web & addrb_valid) 
        ram_cell[addrbl] <= dinb;

endmodule

//����˵��
    //ͬ����дbram��a��ֻ��������ȡָ��b�ڿɶ�д���������debug_module���ж�д
    //дʹ��Ϊ1bit����֧��byte write
//����
    //clk               ����ʱ��
    //addra             a�ڶ���ַ
    //addrb             b�ڶ�д��ַ
    //dinb              b��д��������
    //web               b��дʹ��
//���
    //douta             a�ڶ�����
    //doutb             b�ڶ�����
//ʵ��Ҫ��  
    //�����޸�